library verilog;
use verilog.vl_types.all;
entity checkModule is
end checkModule;
