library verilog;
use verilog.vl_types.all;
entity testBenchAlu is
end testBenchAlu;
