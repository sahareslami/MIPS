library verilog;
use verilog.vl_types.all;
entity testBenchMips is
end testBenchMips;
