library verilog;
use verilog.vl_types.all;
entity testBenchDmem is
end testBenchDmem;
