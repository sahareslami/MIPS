library verilog;
use verilog.vl_types.all;
entity testBenchRegFile is
end testBenchRegFile;
