library verilog;
use verilog.vl_types.all;
entity testBenchIMem is
end testBenchIMem;
