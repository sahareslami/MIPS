library verilog;
use verilog.vl_types.all;
entity TestBenchPc is
end TestBenchPc;
